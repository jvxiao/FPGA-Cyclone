library verilog;
use verilog.vl_types.all;
entity digitalclock_vlg_vec_tst is
end digitalclock_vlg_vec_tst;
