library verilog;
use verilog.vl_types.all;
entity Counter6_vlg_vec_tst is
end Counter6_vlg_vec_tst;
