library verilog;
use verilog.vl_types.all;
entity top_clock_vlg_vec_tst is
end top_clock_vlg_vec_tst;
