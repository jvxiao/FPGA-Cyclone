library verilog;
use verilog.vl_types.all;
entity Quanjia_vlg_check_tst is
    port(
        ci1             : in     vl_logic;
        si              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Quanjia_vlg_check_tst;
