library verilog;
use verilog.vl_types.all;
entity Quanjia_vlg_vec_tst is
end Quanjia_vlg_vec_tst;
