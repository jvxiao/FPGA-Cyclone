module freq(clk,rst_n,clk_1s,clk_1ms,clk_20ms);

input clk,rst_n;

output reg clk_1s,clk_1ms,clk_20ms;

reg [30:0]counter;//1s计数
reg [30:0]cnt1ms;//1ms计数
reg [30:0]cnt;//20ms计数


//1ms
always@(posedge clk or negedge rst_n)
  begin 
	if(!rst_n)
     begin
	    cnt1ms<=0;
       clk_1ms<=0;
     end
   else if(cnt1ms<250)//25000000时间为1s，12500000为0.5s
       cnt1ms<=cnt1ms+1;
	else 
	  begin
       cnt1ms<=0;
		 clk_1ms<=~clk_1ms;
     end
  end


//20ms
always@(posedge clk or negedge rst_n)
  begin 
	if(!rst_n)
     begin
       cnt<=0;
       clk_20ms<=0;
     end
   else if(cnt<50)//25000000时间为1s，12500000为0.5s
       cnt<=cnt+1;
	else 
	  begin
       cnt<=0;
		 clk_20ms<=~clk_20ms;
     end
  end



//1s分频
always@(posedge clk or negedge rst_n)
  begin 
	if(!rst_n)
     begin
       counter<=0;
       clk_1s<=0;
     end
   else if(counter<250)//25000000时间为1s，12500000为0.5s
       counter<=counter+1;
	else 
	  begin
       counter<=0;
		 clk_1s<=~clk_1s;
     end
  end
  
endmodule
