library verilog;
use verilog.vl_types.all;
entity sig_vlg_vec_tst is
end sig_vlg_vec_tst;
